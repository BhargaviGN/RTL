module seq_detector (
    input in, clk, rst, output reg out
);
    
endmodule